LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE hdmi_parameters IS 
    SUBTYPE byte IS STD_LOGIC_VECTOR(7 DOWNTO 0);
    SUBTYPE rgb_t IS STD_LOGIC_VECTOR(23 DOWNTO 0);
    
    CONSTANT FRAME_WIDTH   : INTEGER := 640;
    CONSTANT H_FRONT_PORCH : INTEGER := 16;
    CONSTANT H_BACK_PORCH  : INTEGER := 48;
    CONSTANT H_PULSE_WIDTH : INTEGER := 96;
    CONSTANT H_BLANK       : INTEGER := H_FRONT_PORCH + H_BACK_PORCH + H_PULSE_WIDTH;
    
    CONSTANT FRAME_HEIGHT    : INTEGER := 480;
    CONSTANT V_FRONT_PORCH   : INTEGER := 10;
    CONSTANT V_BACK_PORCH    : INTEGER := 33;
    CONSTANT V_PULSE_WIDTH   : INTEGER := 2;
    CONSTANT V_BLANK         : INTEGER := V_FRONT_PORCH + V_BACK_PORCH + V_PULSE_WIDTH;
    
    CONSTANT H_MAX : INTEGER := FRAME_WIDTH + H_BLANK;
    CONSTANT V_MAX : INTEGER := FRAME_HEIGHT + V_BLANK;
	
	CONSTANT DISPLAY_RESOLUTION : INTEGER := FRAME_WIDTH*FRAME_HEIGHT;
	CONSTANT MAX_RESOLUTION : INTEGER := H_MAX*V_MAX;  

END hdmi_parameters;
